module top();
    reg clk;
    reg reset;
    wire mem_read,mem_write;
    wire [15:0] adr;
    wire [31:0] data;
    wire [31:0] mem_data;

endmodule