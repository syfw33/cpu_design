module controller(
    
);

endmodule